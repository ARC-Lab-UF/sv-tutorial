
// ------SIGNED--------
// 8 bit : byte
// 16 bit: short int
// 32 bit: int
// 64 bit: long int