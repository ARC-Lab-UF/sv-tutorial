// Greg Stitt
// University of Florida

`timescale 1 ns / 100 ps

// Module: moore_tb
// Description: Testbench for the moore module, which implements a Moore FSM.
// Note that if more is changed to use the 1-process version, this testbench
// will start to report errors because of the 1-cycle delay for the outputs.
// It is left as an exercise to adapt the testbench to work for both models.

module moore_tb;

   localparam NUM_CYCLES = 1000;   
   logic clk=0, rst, en;
   logic [3:0] out;

   moore DUT (.*);

   initial begin : generate_clock
      while(1)
	#10 clk = ~clk;      
   end

   logic [$bits(out)-1:0] correct_out;
      
   initial begin
      $timeformat(-9, 0, " ns");

      rst = 1'b1;
      en = 1'b0;
      correct_out = "0001";      
      for (int i=0; i < 5; i++)
	@(posedge clk);

      rst = 1'b0;
      
      for (int i=0; i < NUM_CYCLES; i++) begin
	 en = $random;
	 @(negedge clk);	 
	 if (out != correct_out)
	   $display("ERROR (time %0t): out = %h instead of %h.", $realtime, out, correct_out);
	 @(posedge clk);
	 // The correct output simply rotates every time the enable is asserted.
	 if (en)
	   correct_out = {correct_out[2:0], correct_out[3]};	 	 
      end
            
      disable generate_clock;
      $display("Tests completed.");                    
   end
endmodule
