package accum_tb_pkg;

    localparam int INPUT_WIDTH = 16;    
    localparam int OUTPUT_WIDTH = 32;    

endpackage