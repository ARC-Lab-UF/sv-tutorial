package mult_tb_pkg;

    localparam int INPUT_WIDTH = 16;    

endpackage